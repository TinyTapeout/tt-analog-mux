/// sta-blackbox
(*blackbox*)
module switch_5t(
  input wire en,
  input wire en_b,
  inout wire in,
  inout wire out
);

endmodule // switch_5t