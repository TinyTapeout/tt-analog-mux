VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO switch_5t
  CLASS BLOCK ;
  FOREIGN switch_5t ;
  ORIGIN -0.460 -0.080 ;
  SIZE 14.605 BY 5.560 ;
  PIN VDD
    ANTENNADIFFAREA 5.888800 ;
    PORT
      LAYER nwell ;
        RECT 0.810 2.340 14.885 5.590 ;
      LAYER li1 ;
        RECT 0.990 5.240 14.705 5.410 ;
        RECT 0.990 2.690 1.160 5.240 ;
        RECT 6.930 5.070 8.795 5.240 ;
        RECT 6.930 2.690 7.100 5.070 ;
        RECT 0.990 2.520 7.100 2.690 ;
        RECT 8.595 2.690 8.765 5.070 ;
        RECT 14.535 2.690 14.705 5.240 ;
        RECT 8.595 2.520 14.705 2.690 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 5.394600 ;
    PORT
      LAYER pwell ;
        RECT 0.860 0.080 7.230 2.290 ;
        RECT 8.465 0.080 14.835 2.290 ;
      LAYER li1 ;
        RECT 0.990 1.990 7.100 2.160 ;
        RECT 0.990 0.380 1.160 1.990 ;
        RECT 6.930 0.540 7.100 1.990 ;
        RECT 8.595 1.990 14.705 2.160 ;
        RECT 7.460 1.090 7.630 1.630 ;
        RECT 8.595 0.540 8.765 1.990 ;
        RECT 6.930 0.380 8.765 0.540 ;
        RECT 14.535 0.380 14.705 1.990 ;
        RECT 0.990 0.210 14.705 0.380 ;
        RECT 6.840 0.200 8.830 0.210 ;
      LAYER mcon ;
        RECT 6.930 1.280 7.100 1.450 ;
        RECT 7.460 1.275 7.630 1.445 ;
      LAYER met1 ;
        RECT 6.900 1.615 7.130 1.675 ;
        RECT 6.900 1.610 7.630 1.615 ;
        RECT 6.900 1.115 7.660 1.610 ;
        RECT 6.900 1.055 7.130 1.115 ;
        RECT 7.430 1.110 7.660 1.115 ;
    END
  END VSS
  PIN in
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.040 3.110 2.210 4.510 ;
        RECT 3.000 3.110 3.170 4.510 ;
        RECT 3.960 3.110 4.130 4.510 ;
        RECT 4.920 3.110 5.090 4.510 ;
        RECT 5.880 3.110 6.050 4.510 ;
        RECT 2.040 1.060 2.210 1.620 ;
        RECT 3.000 1.060 3.170 1.620 ;
        RECT 3.960 1.060 4.130 1.620 ;
        RECT 4.920 1.060 5.090 1.620 ;
        RECT 5.880 1.060 6.050 1.620 ;
      LAYER mcon ;
        RECT 2.040 4.085 2.210 4.255 ;
        RECT 2.040 3.725 2.210 3.895 ;
        RECT 2.040 3.365 2.210 3.535 ;
        RECT 3.000 4.085 3.170 4.255 ;
        RECT 3.000 3.725 3.170 3.895 ;
        RECT 3.000 3.365 3.170 3.535 ;
        RECT 3.960 4.085 4.130 4.255 ;
        RECT 3.960 3.725 4.130 3.895 ;
        RECT 3.960 3.365 4.130 3.535 ;
        RECT 4.920 4.085 5.090 4.255 ;
        RECT 4.920 3.725 5.090 3.895 ;
        RECT 4.920 3.365 5.090 3.535 ;
        RECT 5.880 4.085 6.050 4.255 ;
        RECT 5.880 3.725 6.050 3.895 ;
        RECT 5.880 3.365 6.050 3.535 ;
        RECT 2.040 1.255 2.210 1.425 ;
        RECT 3.000 1.255 3.170 1.425 ;
        RECT 3.960 1.255 4.130 1.425 ;
        RECT 4.920 1.255 5.090 1.425 ;
        RECT 5.880 1.255 6.050 1.425 ;
      LAYER met1 ;
        RECT 0.810 5.240 6.050 5.410 ;
        RECT 0.810 2.465 0.980 5.240 ;
        RECT 2.040 4.490 2.210 5.240 ;
        RECT 3.000 4.490 3.170 5.240 ;
        RECT 3.960 4.490 4.130 5.240 ;
        RECT 4.920 4.490 5.090 5.240 ;
        RECT 5.880 4.490 6.050 5.240 ;
        RECT 2.010 3.130 2.240 4.490 ;
        RECT 2.970 3.130 3.200 4.490 ;
        RECT 3.930 3.130 4.160 4.490 ;
        RECT 4.890 3.130 5.120 4.490 ;
        RECT 5.850 3.130 6.080 4.490 ;
        RECT 0.460 2.205 0.980 2.465 ;
        RECT 0.810 0.370 0.980 2.205 ;
        RECT 2.010 1.080 2.240 1.600 ;
        RECT 2.970 1.080 3.200 1.600 ;
        RECT 3.930 1.080 4.160 1.600 ;
        RECT 4.890 1.080 5.120 1.600 ;
        RECT 5.850 1.080 6.080 1.600 ;
        RECT 2.040 0.370 2.210 1.080 ;
        RECT 3.000 0.370 3.170 1.080 ;
        RECT 3.960 0.370 4.130 1.080 ;
        RECT 4.920 0.370 5.090 1.080 ;
        RECT 5.880 0.370 6.050 1.080 ;
        RECT 0.810 0.200 6.050 0.370 ;
    END
  END in
  PIN out
    ANTENNADIFFAREA 3.647200 ;
    PORT
      LAYER li1 ;
        RECT 9.165 3.110 9.335 4.510 ;
        RECT 10.125 3.110 10.295 4.510 ;
        RECT 11.085 3.110 11.255 4.510 ;
        RECT 12.045 3.110 12.215 4.510 ;
        RECT 13.005 3.110 13.175 4.510 ;
        RECT 13.965 3.110 14.135 4.510 ;
        RECT 9.165 1.060 9.335 1.620 ;
        RECT 10.125 1.060 10.295 1.620 ;
        RECT 11.085 1.060 11.255 1.620 ;
        RECT 12.045 1.060 12.215 1.620 ;
        RECT 13.005 1.060 13.175 1.620 ;
        RECT 13.965 1.060 14.135 1.620 ;
      LAYER mcon ;
        RECT 9.165 4.085 9.335 4.255 ;
        RECT 9.165 3.725 9.335 3.895 ;
        RECT 9.165 3.365 9.335 3.535 ;
        RECT 10.125 4.085 10.295 4.255 ;
        RECT 10.125 3.725 10.295 3.895 ;
        RECT 10.125 3.365 10.295 3.535 ;
        RECT 11.085 4.085 11.255 4.255 ;
        RECT 11.085 3.725 11.255 3.895 ;
        RECT 11.085 3.365 11.255 3.535 ;
        RECT 12.045 4.085 12.215 4.255 ;
        RECT 12.045 3.725 12.215 3.895 ;
        RECT 12.045 3.365 12.215 3.535 ;
        RECT 13.005 4.085 13.175 4.255 ;
        RECT 13.005 3.725 13.175 3.895 ;
        RECT 13.005 3.365 13.175 3.535 ;
        RECT 13.965 4.085 14.135 4.255 ;
        RECT 13.965 3.725 14.135 3.895 ;
        RECT 13.965 3.365 14.135 3.535 ;
        RECT 9.165 1.255 9.335 1.425 ;
        RECT 10.125 1.255 10.295 1.425 ;
        RECT 11.085 1.255 11.255 1.425 ;
        RECT 12.045 1.255 12.215 1.425 ;
        RECT 13.005 1.255 13.175 1.425 ;
        RECT 13.965 1.255 14.135 1.425 ;
      LAYER met1 ;
        RECT 9.135 3.130 9.365 4.490 ;
        RECT 10.095 3.130 10.325 4.490 ;
        RECT 11.055 3.130 11.285 4.490 ;
        RECT 12.015 3.130 12.245 4.490 ;
        RECT 12.975 3.130 13.205 4.490 ;
        RECT 13.935 3.130 14.165 4.490 ;
        RECT 9.165 2.425 9.335 3.130 ;
        RECT 10.125 2.425 10.295 3.130 ;
        RECT 11.085 2.425 11.255 3.130 ;
        RECT 12.045 2.425 12.215 3.130 ;
        RECT 13.005 2.425 13.175 3.130 ;
        RECT 13.965 2.425 14.135 3.130 ;
        RECT 9.165 2.255 14.710 2.425 ;
        RECT 9.165 1.600 9.335 2.255 ;
        RECT 10.125 1.600 10.295 2.255 ;
        RECT 11.085 1.600 11.255 2.255 ;
        RECT 12.045 1.600 12.215 2.255 ;
        RECT 13.005 1.600 13.175 2.255 ;
        RECT 13.965 1.600 14.135 2.255 ;
        RECT 9.135 1.080 9.365 1.600 ;
        RECT 10.095 1.080 10.325 1.600 ;
        RECT 11.055 1.080 11.285 1.600 ;
        RECT 12.015 1.080 12.245 1.600 ;
        RECT 12.975 1.080 13.205 1.600 ;
        RECT 13.935 1.080 14.165 1.600 ;
    END
  END out
  PIN en
    ANTENNAGATEAREA 1.560000 ;
    PORT
      LAYER li1 ;
        RECT 1.480 0.635 6.610 0.885 ;
        RECT 9.085 0.635 14.215 0.885 ;
      LAYER mcon ;
        RECT 1.560 0.675 1.730 0.845 ;
        RECT 6.360 0.675 6.530 0.845 ;
        RECT 9.165 0.675 9.335 0.845 ;
        RECT 13.965 0.675 14.135 0.845 ;
      LAYER met1 ;
        RECT 1.460 0.620 1.820 0.880 ;
        RECT 6.270 0.630 6.630 0.890 ;
        RECT 9.075 0.630 9.435 0.890 ;
        RECT 13.875 0.630 14.235 0.890 ;
      LAYER via ;
        RECT 1.510 0.620 1.770 0.880 ;
        RECT 6.320 0.630 6.580 0.890 ;
        RECT 9.125 0.630 9.385 0.890 ;
        RECT 13.925 0.630 14.185 0.890 ;
      LAYER met2 ;
        RECT 1.510 0.915 1.770 0.930 ;
        RECT 1.970 0.915 2.300 0.925 ;
        RECT 6.320 0.915 6.580 0.940 ;
        RECT 9.125 0.915 9.385 0.940 ;
        RECT 13.925 0.915 14.185 0.940 ;
        RECT 0.460 0.655 14.185 0.915 ;
        RECT 1.510 0.570 1.770 0.655 ;
        RECT 1.970 0.595 2.300 0.655 ;
        RECT 6.320 0.580 6.580 0.655 ;
        RECT 9.125 0.580 9.385 0.655 ;
        RECT 13.925 0.580 14.185 0.655 ;
    END
  END en
  PIN en_b
    ANTENNAGATEAREA 4.155000 ;
    PORT
      LAYER li1 ;
        RECT 1.480 4.690 6.610 4.940 ;
        RECT 9.085 4.690 14.215 4.940 ;
        RECT 7.600 1.800 7.930 1.970 ;
      LAYER mcon ;
        RECT 1.560 4.730 1.730 4.900 ;
        RECT 6.360 4.730 6.530 4.900 ;
        RECT 9.165 4.730 9.335 4.900 ;
        RECT 13.965 4.730 14.135 4.900 ;
        RECT 7.680 1.800 7.850 1.970 ;
      LAYER met1 ;
        RECT 1.465 4.685 1.825 4.945 ;
        RECT 6.260 4.690 6.620 4.950 ;
        RECT 9.065 4.690 9.425 4.950 ;
        RECT 13.865 4.690 14.225 4.950 ;
        RECT 7.585 1.805 7.945 2.065 ;
        RECT 7.620 1.770 7.910 1.805 ;
      LAYER via ;
        RECT 1.515 4.685 1.775 4.945 ;
        RECT 6.310 4.690 6.570 4.950 ;
        RECT 9.115 4.690 9.375 4.950 ;
        RECT 13.915 4.690 14.175 4.950 ;
        RECT 7.635 1.805 7.895 2.065 ;
      LAYER met2 ;
        RECT 1.515 4.950 1.775 4.995 ;
        RECT 6.310 4.950 6.570 5.000 ;
        RECT 9.115 4.950 9.375 5.000 ;
        RECT 13.915 4.950 14.175 5.000 ;
        RECT 0.505 4.690 14.245 4.950 ;
        RECT 1.515 4.635 1.775 4.690 ;
        RECT 6.310 4.640 6.570 4.690 ;
        RECT 7.635 1.755 7.895 4.690 ;
        RECT 9.115 4.640 9.375 4.690 ;
        RECT 13.915 4.640 14.175 4.690 ;
    END
  END en_b
  OBS
      LAYER pwell ;
        RECT 7.270 0.980 8.260 1.740 ;
      LAYER li1 ;
        RECT 1.560 3.110 1.730 4.510 ;
        RECT 2.520 3.110 2.690 4.510 ;
        RECT 3.480 3.110 3.650 4.510 ;
        RECT 4.440 3.110 4.610 4.510 ;
        RECT 5.400 3.110 5.570 4.510 ;
        RECT 6.360 3.110 6.530 4.510 ;
        RECT 9.645 3.110 9.815 4.510 ;
        RECT 10.605 3.110 10.775 4.510 ;
        RECT 11.565 3.110 11.735 4.510 ;
        RECT 12.525 3.110 12.695 4.510 ;
        RECT 13.485 3.110 13.655 4.510 ;
        RECT 1.560 1.060 1.730 1.620 ;
        RECT 2.520 1.060 2.690 1.620 ;
        RECT 3.480 1.060 3.650 1.620 ;
        RECT 4.440 1.060 4.610 1.620 ;
        RECT 5.400 1.060 5.570 1.620 ;
        RECT 6.360 1.060 6.530 1.620 ;
        RECT 7.900 1.090 8.070 1.630 ;
        RECT 9.645 1.060 9.815 1.620 ;
        RECT 10.605 1.060 10.775 1.620 ;
        RECT 11.565 1.060 11.735 1.620 ;
        RECT 12.525 1.060 12.695 1.620 ;
        RECT 13.485 1.060 13.655 1.620 ;
      LAYER mcon ;
        RECT 1.560 4.085 1.730 4.255 ;
        RECT 1.560 3.725 1.730 3.895 ;
        RECT 1.560 3.365 1.730 3.535 ;
        RECT 2.520 4.085 2.690 4.255 ;
        RECT 2.520 3.725 2.690 3.895 ;
        RECT 2.520 3.365 2.690 3.535 ;
        RECT 3.480 4.085 3.650 4.255 ;
        RECT 3.480 3.725 3.650 3.895 ;
        RECT 3.480 3.365 3.650 3.535 ;
        RECT 4.440 4.085 4.610 4.255 ;
        RECT 4.440 3.725 4.610 3.895 ;
        RECT 4.440 3.365 4.610 3.535 ;
        RECT 5.400 4.085 5.570 4.255 ;
        RECT 5.400 3.725 5.570 3.895 ;
        RECT 5.400 3.365 5.570 3.535 ;
        RECT 6.360 4.085 6.530 4.255 ;
        RECT 6.360 3.725 6.530 3.895 ;
        RECT 6.360 3.365 6.530 3.535 ;
        RECT 9.645 4.085 9.815 4.255 ;
        RECT 9.645 3.725 9.815 3.895 ;
        RECT 9.645 3.365 9.815 3.535 ;
        RECT 10.605 4.085 10.775 4.255 ;
        RECT 10.605 3.725 10.775 3.895 ;
        RECT 10.605 3.365 10.775 3.535 ;
        RECT 11.565 4.085 11.735 4.255 ;
        RECT 11.565 3.725 11.735 3.895 ;
        RECT 11.565 3.365 11.735 3.535 ;
        RECT 12.525 4.085 12.695 4.255 ;
        RECT 12.525 3.725 12.695 3.895 ;
        RECT 12.525 3.365 12.695 3.535 ;
        RECT 13.485 4.085 13.655 4.255 ;
        RECT 13.485 3.725 13.655 3.895 ;
        RECT 13.485 3.365 13.655 3.535 ;
        RECT 1.560 1.255 1.730 1.425 ;
        RECT 2.520 1.255 2.690 1.425 ;
        RECT 3.480 1.255 3.650 1.425 ;
        RECT 4.440 1.255 4.610 1.425 ;
        RECT 5.400 1.255 5.570 1.425 ;
        RECT 6.360 1.255 6.530 1.425 ;
        RECT 7.900 1.275 8.070 1.445 ;
        RECT 9.645 1.255 9.815 1.425 ;
        RECT 10.605 1.255 10.775 1.425 ;
        RECT 11.565 1.255 11.735 1.425 ;
        RECT 12.525 1.255 12.695 1.425 ;
        RECT 13.485 1.255 13.655 1.425 ;
      LAYER met1 ;
        RECT 8.415 5.240 13.655 5.410 ;
        RECT 1.530 3.130 1.760 4.490 ;
        RECT 2.490 3.130 2.720 4.490 ;
        RECT 3.450 3.130 3.680 4.490 ;
        RECT 4.410 3.130 4.640 4.490 ;
        RECT 5.370 3.130 5.600 4.490 ;
        RECT 6.330 3.130 6.560 4.490 ;
        RECT 1.560 2.425 1.730 3.130 ;
        RECT 2.520 2.425 2.690 3.130 ;
        RECT 3.480 2.425 3.650 3.130 ;
        RECT 4.440 2.425 4.610 3.130 ;
        RECT 5.400 2.425 5.570 3.130 ;
        RECT 6.360 2.425 6.530 3.130 ;
        RECT 8.415 2.425 8.585 5.240 ;
        RECT 9.645 4.490 9.815 5.240 ;
        RECT 10.605 4.490 10.775 5.240 ;
        RECT 11.565 4.490 11.735 5.240 ;
        RECT 12.525 4.490 12.695 5.240 ;
        RECT 13.485 4.490 13.655 5.240 ;
        RECT 9.615 3.130 9.845 4.490 ;
        RECT 10.575 3.130 10.805 4.490 ;
        RECT 11.535 3.130 11.765 4.490 ;
        RECT 12.495 3.130 12.725 4.490 ;
        RECT 13.455 3.130 13.685 4.490 ;
        RECT 1.560 2.255 8.585 2.425 ;
        RECT 1.560 1.600 1.730 2.255 ;
        RECT 2.520 1.600 2.690 2.255 ;
        RECT 3.480 1.600 3.650 2.255 ;
        RECT 4.440 1.600 4.610 2.255 ;
        RECT 5.400 1.600 5.570 2.255 ;
        RECT 6.360 1.600 6.530 2.255 ;
        RECT 8.415 1.615 8.585 2.255 ;
        RECT 7.900 1.610 8.585 1.615 ;
        RECT 1.530 1.080 1.760 1.600 ;
        RECT 2.490 1.080 2.720 1.600 ;
        RECT 3.450 1.080 3.680 1.600 ;
        RECT 4.410 1.080 4.640 1.600 ;
        RECT 5.370 1.080 5.600 1.600 ;
        RECT 6.330 1.080 6.560 1.600 ;
        RECT 7.870 1.115 8.585 1.610 ;
        RECT 7.870 1.110 8.100 1.115 ;
        RECT 8.415 0.370 8.585 1.115 ;
        RECT 9.615 1.080 9.845 1.600 ;
        RECT 10.575 1.080 10.805 1.600 ;
        RECT 11.535 1.080 11.765 1.600 ;
        RECT 12.495 1.080 12.725 1.600 ;
        RECT 13.455 1.080 13.685 1.600 ;
        RECT 9.645 0.370 9.815 1.080 ;
        RECT 10.605 0.370 10.775 1.080 ;
        RECT 11.565 0.370 11.735 1.080 ;
        RECT 12.525 0.370 12.695 1.080 ;
        RECT 13.485 0.370 13.655 1.080 ;
        RECT 8.415 0.200 13.655 0.370 ;
  END
END switch_5t
END LIBRARY

